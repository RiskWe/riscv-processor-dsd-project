`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:15:33 10/10/2024 
// Design Name: 
// Module Name:    AND_logic 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module AND_logic(branch, zero, and_out);

input branch, zero;
output and_out;
output and_out;

assign and_out = branch & zero;
endmodule
