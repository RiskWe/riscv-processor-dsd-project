`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:36:30 10/09/2024 
// Design Name: 
// Module Name:    PC 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module PC(clk, reset, PC_in, PC_out);

input clk, reset;
input 	 [31:0] PC_in;
input reg [31:0] PC_out;

always @(posedge clk or posedge reset)
begin
if(reset)
	PC_out <= 32'b00;
else
	PC_out <= PC_in;
end

endmodule
